

`include "uvm_macros.svh"
package axi4_sram_tests_pkg;
	import uvm_pkg::*;
	import axi4_sram_env_pkg::*;
	import Axi4SramTestsBasePkg::*;
	
	`include "axi4_sram_test_base.svh"
	
endpackage
