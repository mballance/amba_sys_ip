/****************************************************************************
 * Axi4SramTestsBasePkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: Axi4SramTestsBasePkg
 * 
 * TODO: Add package documentation
 */
package Axi4SramTestsBasePkg;
	import uvm_pkg::*;

	`include "Axi4SramTestBase.svh"

endpackage


