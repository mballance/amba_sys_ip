/****************************************************************************
 * Axi4SramEnvBasePkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: Axi4SramEnvBasePkg
 * 
 * TODO: Add package documentation
 */
package Axi4SramEnvBasePkg;
	import uvm_pkg::*;

	`include "Axi4SramEnvBase.svh"

endpackage


