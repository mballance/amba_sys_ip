
`include "uvm_macros.svh"

package axi4_sram_env_pkg;
	import uvm_pkg::*;
	import Axi4SramEnvBasePkg::*;

	`include "axi4_sram_env.svh"
	
endpackage
